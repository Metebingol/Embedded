library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity JA_pin_manager_v1_0_S00_AXI is
	generic (
		-- Users to add parameters here
        outType1                 : string := "StandardIO"; -- "PWM" and "PULSE"
        outType2                 : string := "StandardIO"; -- "PWM" and "PULSE"
        outType3                 : string := "StandardIO"; -- "PWM" and "PULSE"
        outType4                 : string := "StandardIO"; -- "PWM" and "PULSE"
        outType5                 : string := "StandardIO"; -- "PWM" and "PULSE"
        outType6                 : string := "StandardIO"; -- "PWM" and "PULSE"
        outType7                 : string := "StandardIO"; -- "PWM" and "PULSE"
        outType8                 : string := "StandardIO"; -- "PWM" and "PULSE"
        pwmFrequency1            : integer := 20;
        pwmFrequency2            : integer := 20;
        pwmFrequency3            : integer := 20;
        pwmFrequency4            : integer := 20;
        pwmFrequency5            : integer := 20;
        pwmFrequency6            : integer := 20;
        pwmFrequency7            : integer := 20;
        pwmFrequency8            : integer := 20;
		-- User parameters ends
		-- Do not modify the parameters beyond this line

		-- Width of S_AXI data bus
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		-- Width of S_AXI address bus
		C_S_AXI_ADDR_WIDTH	: integer	:= 4
	);
	port (
		-- Users to add ports here
        JAoutputPin1            : inout std_logic := '0';
        JAoutputPin2            : inout std_logic := '0';
        JAoutputPin3            : inout std_logic := '0';
        JAoutputPin4            : inout std_logic := '0';
        JAoutputPin5            : inout std_logic := '0';
        JAoutputPin6            : inout std_logic := '0';
        JAoutputPin7            : inout std_logic := '0';
        JAoutputPin8            : inout std_logic := '0';
		-- User ports ends
		-- Do not modify the ports beyond this line

		-- Global Clock Signal
		S_AXI_ACLK	: in std_logic;
		-- Global Reset Signal. This Signal is Active LOW
		S_AXI_ARESETN	: in std_logic;
		-- Write address (issued by master, acceped by Slave)
		S_AXI_AWADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		-- Write channel Protection type. This signal indicates the
    		-- privilege and security level of the transaction, and whether
    		-- the transaction is a data access or an instruction access.
		S_AXI_AWPROT	: in std_logic_vector(2 downto 0);
		-- Write address valid. This signal indicates that the master signaling
    		-- valid write address and control information.
		S_AXI_AWVALID	: in std_logic;
		-- Write address ready. This signal indicates that the slave is ready
    		-- to accept an address and associated control signals.
		S_AXI_AWREADY	: out std_logic;
		-- Write data (issued by master, acceped by Slave) 
		S_AXI_WDATA	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		-- Write strobes. This signal indicates which byte lanes hold
    		-- valid data. There is one write strobe bit for each eight
    		-- bits of the write data bus.    
		S_AXI_WSTRB	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		-- Write valid. This signal indicates that valid write
    		-- data and strobes are available.
		S_AXI_WVALID	: in std_logic;
		-- Write ready. This signal indicates that the slave
    		-- can accept the write data.
		S_AXI_WREADY	: out std_logic;
		-- Write response. This signal indicates the status
    		-- of the write transaction.
		S_AXI_BRESP	: out std_logic_vector(1 downto 0);
		-- Write response valid. This signal indicates that the channel
    		-- is signaling a valid write response.
		S_AXI_BVALID	: out std_logic;
		-- Response ready. This signal indicates that the master
    		-- can accept a write response.
		S_AXI_BREADY	: in std_logic;
		-- Read address (issued by master, acceped by Slave)
		S_AXI_ARADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		-- Protection type. This signal indicates the privilege
    		-- and security level of the transaction, and whether the
    		-- transaction is a data access or an instruction access.
		S_AXI_ARPROT	: in std_logic_vector(2 downto 0);
		-- Read address valid. This signal indicates that the channel
    		-- is signaling valid read address and control information.
		S_AXI_ARVALID	: in std_logic;
		-- Read address ready. This signal indicates that the slave is
    		-- ready to accept an address and associated control signals.
		S_AXI_ARREADY	: out std_logic;
		-- Read data (issued by slave)
		S_AXI_RDATA	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		-- Read response. This signal indicates the status of the
    		-- read transfer.
		S_AXI_RRESP	: out std_logic_vector(1 downto 0);
		-- Read valid. This signal indicates that the channel is
    		-- signaling the required read data.
		S_AXI_RVALID	: out std_logic;
		-- Read ready. This signal indicates that the master can
    		-- accept the read data and response information.
		S_AXI_RREADY	: in std_logic
	);
end JA_pin_manager_v1_0_S00_AXI;

architecture arch_imp of JA_pin_manager_v1_0_S00_AXI is

	-- AXI4LITE signals
	signal axi_awaddr	: std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
	signal axi_awready	: std_logic;
	signal axi_wready	: std_logic;
	signal axi_bresp	: std_logic_vector(1 downto 0);
	signal axi_bvalid	: std_logic;
	signal axi_araddr	: std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
	signal axi_arready	: std_logic;
	signal axi_rdata	: std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal axi_rresp	: std_logic_vector(1 downto 0);
	signal axi_rvalid	: std_logic;

	-- Example-specific design signals
	-- local parameter for addressing 32 bit / 64 bit C_S_AXI_DATA_WIDTH
	-- ADDR_LSB is used for addressing 32/64 bit registers/memories
	-- ADDR_LSB = 2 for 32 bits (n downto 2)
	-- ADDR_LSB = 3 for 64 bits (n downto 3)
	constant ADDR_LSB  : integer := (C_S_AXI_DATA_WIDTH/32)+ 1;
	constant OPT_MEM_ADDR_BITS : integer := 1;
	------------------------------------------------
	---- Signals for user logic register space example
	--------------------------------------------------
	---- Number of Slave Registers 4
	signal slv_reg0	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0); -- enable (8bit) Output Standard (8bit) 
	signal slv_reg1	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0); -- pwm percent 
	signal slv_reg2	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0); -- pulse number 
	signal slv_reg3	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0); -- busy(8bit) -- type(16bit) example: "11111111-00000000-11,11,11,11,11,11,11,11 (11:IOStandard 10:PWM 01:pulse 00:NW)"
	signal slv_reg_rden	: std_logic;
	signal slv_reg_wren	: std_logic;
	signal reg_data_out	:std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal byte_index	: integer;
	signal aw_en	: std_logic;

begin
	-- I/O Connections assignments

	S_AXI_AWREADY	<= axi_awready;
	S_AXI_WREADY	<= axi_wready;
	S_AXI_BRESP	<= axi_bresp;
	S_AXI_BVALID	<= axi_bvalid;
	S_AXI_ARREADY	<= axi_arready;
	S_AXI_RDATA	<= axi_rdata;
	S_AXI_RRESP	<= axi_rresp;
	S_AXI_RVALID	<= axi_rvalid;
	-- Implement axi_awready generation
	-- axi_awready is asserted for one S_AXI_ACLK clock cycle when both
	-- S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_awready is
	-- de-asserted when reset is low.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_awready <= '0';
	      aw_en <= '1';
	    else
	      if (axi_awready = '0' and S_AXI_AWVALID = '1' and S_AXI_WVALID = '1' and aw_en = '1') then
	        -- slave is ready to accept write address when
	        -- there is a valid write address and write data
	        -- on the write address and data bus. This design 
	        -- expects no outstanding transactions. 
	           axi_awready <= '1';
	           aw_en <= '0';
	        elsif (S_AXI_BREADY = '1' and axi_bvalid = '1') then
	           aw_en <= '1';
	           axi_awready <= '0';
	      else
	        axi_awready <= '0';
	      end if;
	    end if;
	  end if;
	end process;

	-- Implement axi_awaddr latching
	-- This process is used to latch the address when both 
	-- S_AXI_AWVALID and S_AXI_WVALID are valid. 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_awaddr <= (others => '0');
	    else
	      if (axi_awready = '0' and S_AXI_AWVALID = '1' and S_AXI_WVALID = '1' and aw_en = '1') then
	        -- Write Address latching
	        axi_awaddr <= S_AXI_AWADDR;
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement axi_wready generation
	-- axi_wready is asserted for one S_AXI_ACLK clock cycle when both
	-- S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_wready is 
	-- de-asserted when reset is low. 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_wready <= '0';
	    else
	      if (axi_wready = '0' and S_AXI_WVALID = '1' and S_AXI_AWVALID = '1' and aw_en = '1') then
	          -- slave is ready to accept write data when 
	          -- there is a valid write address and write data
	          -- on the write address and data bus. This design 
	          -- expects no outstanding transactions.           
	          axi_wready <= '1';
	      else
	        axi_wready <= '0';
	      end if;
	    end if;
	  end if;
	end process; 

	-- Implement memory mapped register select and write logic generation
	-- The write data is accepted and written to memory mapped registers when
	-- axi_awready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted. Write strobes are used to
	-- select byte enables of slave registers while writing.
	-- These registers are cleared when reset (active low) is applied.
	-- Slave register write enable is asserted when valid address and data are available
	-- and the slave is ready to accept the write address and write data.
	slv_reg_wren <= axi_wready and S_AXI_WVALID and axi_awready and S_AXI_AWVALID ;

	process (S_AXI_ACLK)
	variable loc_addr :std_logic_vector(OPT_MEM_ADDR_BITS downto 0); 
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      slv_reg0 <= (others => '0');
	      slv_reg1 <= (others => '0');
	      slv_reg2 <= (others => '0');
	      slv_reg3 <= (others => '0');
	    else
	      loc_addr := axi_awaddr(ADDR_LSB + OPT_MEM_ADDR_BITS downto ADDR_LSB);
	      if (slv_reg_wren = '1') then
	        case loc_addr is
	          when b"00" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 0
	                slv_reg0(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 1
	                slv_reg1(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 2
	                slv_reg2(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"11" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 3
	                slv_reg3(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when others =>
	            slv_reg0 <= slv_reg0;
	            slv_reg1 <= slv_reg1;
	            slv_reg2 <= slv_reg2;
	            slv_reg3 <= slv_reg3;
	        end case;
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement write response logic generation
	-- The write response and response valid signals are asserted by the slave 
	-- when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.  
	-- This marks the acceptance of address and indicates the status of 
	-- write transaction.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_bvalid  <= '0';
	      axi_bresp   <= "00"; --need to work more on the responses
	    else
	      if (axi_awready = '1' and S_AXI_AWVALID = '1' and axi_wready = '1' and S_AXI_WVALID = '1' and axi_bvalid = '0'  ) then
	        axi_bvalid <= '1';
	        axi_bresp  <= "00"; 
	      elsif (S_AXI_BREADY = '1' and axi_bvalid = '1') then   --check if bready is asserted while bvalid is high)
	        axi_bvalid <= '0';                                 -- (there is a possibility that bready is always asserted high)
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement axi_arready generation
	-- axi_arready is asserted for one S_AXI_ACLK clock cycle when
	-- S_AXI_ARVALID is asserted. axi_awready is 
	-- de-asserted when reset (active low) is asserted. 
	-- The read address is also latched when S_AXI_ARVALID is 
	-- asserted. axi_araddr is reset to zero on reset assertion.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_arready <= '0';
	      axi_araddr  <= (others => '1');
	    else
	      if (axi_arready = '0' and S_AXI_ARVALID = '1') then
	        -- indicates that the slave has acceped the valid read address
	        axi_arready <= '1';
	        -- Read Address latching 
	        axi_araddr  <= S_AXI_ARADDR;           
	      else
	        axi_arready <= '0';
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement axi_arvalid generation
	-- axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both 
	-- S_AXI_ARVALID and axi_arready are asserted. The slave registers 
	-- data are available on the axi_rdata bus at this instance. The 
	-- assertion of axi_rvalid marks the validity of read data on the 
	-- bus and axi_rresp indicates the status of read transaction.axi_rvalid 
	-- is deasserted on reset (active low). axi_rresp and axi_rdata are 
	-- cleared to zero on reset (active low).  
	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then
	    if S_AXI_ARESETN = '0' then
	      axi_rvalid <= '0';
	      axi_rresp  <= "00";
	    else
	      if (axi_arready = '1' and S_AXI_ARVALID = '1' and axi_rvalid = '0') then
	        -- Valid read data is available at the read data bus
	        axi_rvalid <= '1';
	        axi_rresp  <= "00"; -- 'OKAY' response
	      elsif (axi_rvalid = '1' and S_AXI_RREADY = '1') then
	        -- Read data is accepted by the master
	        axi_rvalid <= '0';
	      end if;            
	    end if;
	  end if;
	end process;

	-- Implement memory mapped register select and read logic generation
	-- Slave register read enable is asserted when valid address is available
	-- and the slave is ready to accept the read address.
	slv_reg_rden <= axi_arready and S_AXI_ARVALID and (not axi_rvalid) ;

	process (slv_reg0, slv_reg1, slv_reg2, slv_reg3, axi_araddr, S_AXI_ARESETN, slv_reg_rden)
	variable loc_addr :std_logic_vector(OPT_MEM_ADDR_BITS downto 0);
	begin
	    -- Address decoding for reading registers
	    loc_addr := axi_araddr(ADDR_LSB + OPT_MEM_ADDR_BITS downto ADDR_LSB);
	    case loc_addr is
	      when b"00" =>
	        reg_data_out <= slv_reg0;
	      when b"01" =>
	        reg_data_out <= slv_reg1;
	      when b"10" =>
	        reg_data_out <= slv_reg2;
	      when b"11" =>
	        reg_data_out <= slv_reg3;
	      when others =>
	        reg_data_out  <= (others => '0');
	    end case;
	end process; 

	-- Output register or memory read data
	process( S_AXI_ACLK ) is
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	      axi_rdata  <= (others => '0');
	    else
	      if (slv_reg_rden = '1') then
	        -- When there is a valid read address (S_AXI_ARVALID) with 
	        -- acceptance of read address by the slave (axi_arready), 
	        -- output the read dada 
	        -- Read address mux
	          axi_rdata <= reg_data_out;     -- register read data
	      end if;   
	    end if;
	  end if;
	end process;

    

	-- Add user logic here
	-- JA 1 
	process( S_AXI_ACLK ) is
	variable pwmPercent    : integer := 0;
	variable pwmCount      : integer := 100_000_000/(pwmFrequency1*1000);
	variable count         : integer := 0;
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	       axi_rdata  <= (others => '0');
	    else
	       if slv_reg0(0) = '1' then   -- enable for JA1
	           slv_reg3(0) <= '1';     -- busy for JA1
	           case outType1 is 
	               when "StandardIO"   => 
	                   slv_reg3(9 downto 8) <= "11";       -- MODE
	                   if slv_reg_rden = '1' then
	                       JAoutputPin1 <= slv_reg0(8);    -- JA PIN-1 
	                   end if;
	               when "PWM"          => 
	                   slv_reg3(9 downto 8) <= "10";
	                   if slv_reg_rden = '1' then
                           if count >= pwmCount then
                                pwmPercent := to_integer(unsigned(slv_reg1(3 downto 0)));
                                pwmCount := 100_000_000/(pwmFrequency1*1000);
                                count := 0;
                           elsif (count <= (pwmCount*pwmPercent/16)) then
                               JAoutputPin1 <= '1';
                           elsif (count > (pwmCount*pwmPercent/16) and (count < (pwmCount))) then
                               JAoutputPin1 <= '0';
                           end if;
	                   end if;
	                   count := count + 1;
	               when "PULSE"        =>
	                   slv_reg3(9 downto 8) <= "01";
	                   if slv_reg_rden = '1' then
	                       if count = 0 then
	                           count := to_integer(unsigned(slv_reg2(3 downto 0)));
	                       end if;
	                       if count > 2 then
	                           JAoutputPin1 <= not JAoutputPin1;
	                       end if;
	                   end if;
	                   if count > 1 then
	                      count := count -1;
	                   end if;
	               when others         =>
	                   slv_reg3(9 downto 8) <= "00";    
	           end case;
	       else 
	           slv_reg3(0) <= '0'; -- busy for JA1
	           count := 0;
	       end if;
	    end if;
	  end if;
	end process;   
	

	-- JA 2 
	process( S_AXI_ACLK ) is
	variable pwmPercent    : integer := 0;
	variable pwmCount      : integer := 100_000_000/(pwmFrequency2*1000);
	variable count         : integer := 0;
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	       axi_rdata  <= (others => '0');
	    else
	       if slv_reg0(1) = '1' then       -- enable fpr JA2
	           slv_reg3(1) <= '1';         -- busy for JA2
	           case outType2 is 
	               when "StandardIO"   => 
	                   slv_reg3(11 downto 10) <= "11"; -- Mode
	                   if slv_reg_rden = '1' then
	                       JAoutputPin2 <= slv_reg0(9);
	                   end if;
	               when "PWM"          => 
	                   slv_reg3(11 downto 10) <= "10";
	                   if slv_reg_rden = '1' then
                           if count >= pwmCount then
                                pwmPercent := to_integer(unsigned(slv_reg1(7 downto 4)));
                                pwmCount := 100_000_000/(pwmFrequency2*1000);
                                count := 0;
                           elsif (count <= (pwmCount*pwmPercent/16)) then
                               JAoutputPin2 <= '1';
                           elsif (count > (pwmCount*pwmPercent/16) and (count < (pwmCount))) then
                               JAoutputPin2 <= '0';
                           end if;
	                   end if;
	                   count := count + 1;
	               when "PULSE"        =>
	                   slv_reg3(11 downto 10) <= "01";
	                   if slv_reg_rden = '1' then
	                       if count = 0 then
	                           count := to_integer(unsigned(slv_reg2(7 downto 4)));
	                       end if;
	                       if count > 2 then
	                           JAoutputPin2 <= not JAoutputPin2;
	                       end if;
	                   end if;
	                   if count > 1 then
	                      count := count -1;
	                   end if;
	               when others         =>
	                   slv_reg3(11 downto 10) <= "00";    
	           end case;
	       else 
	           slv_reg3(1) <= '0'; -- busy for JA2
	           count := 0;
	       end if;
	    end if;
	  end if;
	end process;   



	-- JA 3
	process( S_AXI_ACLK ) is
	variable pwmPercent    : integer := 0;
	variable pwmCount      : integer := 100_000_000/(pwmFrequency3*1000);
	variable count         : integer := 0;
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	       axi_rdata  <= (others => '0');
	    else
	       if slv_reg0(2) = '1' then   -- enable for JA3
	           slv_reg3(2) <= '1';     -- busy for JA3
	           case outType3 is 
	               when "StandardIO"   => 
	                   slv_reg3(13 downto 12) <= "11";
	                   if slv_reg_rden = '1' then
	                       JAoutputPin3 <= slv_reg0(10);
	                   end if;
	               when "PWM"          => 
	                   slv_reg3(13 downto 12) <= "10";
	                   if slv_reg_rden = '1' then
                           if count >= pwmCount then
                                pwmPercent := to_integer(unsigned(slv_reg1(11 downto 8)));
                                pwmCount := 100_000_000/(pwmFrequency3*1000);
                                count := 0;
                           elsif (count <= (pwmCount*pwmPercent/16)) then
                               JAoutputPin3 <= '1';
                           elsif (count > (pwmCount*pwmPercent/16) and (count < (pwmCount))) then
                               JAoutputPin3 <= '0';
                           end if;
	                   end if;
	                   count := count + 1;
	               when "PULSE"        =>
	                   slv_reg3(13 downto 12) <= "01";
	                   if slv_reg_rden = '1' then
	                       if count = 0 then
	                           count := to_integer(unsigned(slv_reg2(11 downto 8)));
	                       end if;
	                       if count > 2 then
	                           JAoutputPin3 <= not JAoutputPin3;
	                       end if;
	                   end if;
	                   if count > 1 then
	                      count := count -1;
	                   end if;
	               when others         =>
	                   slv_reg3(13 downto 12) <= "00";    
	           end case;
	       else 
	           slv_reg3(2) <= '0'; -- busy for JA3
	           count := 0;
	       end if;
	    end if;
	  end if;
	end process;   



	-- JA 4
	process( S_AXI_ACLK ) is
	variable pwmPercent    : integer := 0;
	variable pwmCount      : integer := 100_000_000/(pwmFrequency4*1000);
	variable count         : integer := 0;
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	       axi_rdata  <= (others => '0');
	    else
	       if slv_reg0(3) = '1' then   -- enable for JA4
	           slv_reg3(3) <= '1';     -- busy for JA4
	           case outType4 is 
	               when "StandardIO"   => 
	                   slv_reg3(15 downto 14) <= "11";
	                   if slv_reg_rden = '1' then
	                       JAoutputPin4 <= slv_reg0(11);
	                   end if;
	               when "PWM"          => 
	                   slv_reg3(15 downto 14) <= "10";
	                   if slv_reg_rden = '1' then
                           if count >= pwmCount then
                                pwmPercent := to_integer(unsigned(slv_reg1(15 downto 12)));
                                pwmCount := 100_000_000/(pwmFrequency4*1000);
                                count := 0;
                           elsif (count <= (pwmCount*pwmPercent/16)) then
                               JAoutputPin4 <= '1';
                           elsif (count > (pwmCount*pwmPercent/16) and (count < (pwmCount))) then
                               JAoutputPin4 <= '0';
                           end if;
	                   end if;
	                   count := count + 1;
	               when "PULSE"        =>
	                   slv_reg3(15 downto 14) <= "01";
	                   if slv_reg_rden = '1' then
	                       if count = 0 then
	                           count := to_integer(unsigned(slv_reg2(15 downto 12)));
	                       end if;
	                       if count > 2 then
	                           JAoutputPin4 <= not JAoutputPin4;
	                       end if;
	                   end if;
	                   if count > 1 then
	                      count := count -1;
	                   end if;
	               when others         =>
	                   slv_reg3(15 downto 14) <= "00";    
	           end case;
	       else 
	           slv_reg3(3) <= '0'; -- busy for JA4
	           count := 0;
	       end if;
	    end if;
	  end if;
	end process;   



	-- JA 5
	process( S_AXI_ACLK ) is
	variable pwmPercent    : integer := 0;
	variable pwmCount      : integer := 100_000_000/(pwmFrequency5*1000);
	variable count         : integer := 0;
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	       axi_rdata  <= (others => '0');
	    else
	       if slv_reg0(4) = '1' then   -- enable for JA5
	           slv_reg3(4) <= '1';     -- busy for JA5
	           case outType5 is 
	               when "StandardIO"   => 
	                   slv_reg3(17 downto 16) <= "11";
	                   if slv_reg_rden = '1' then
	                       JAoutputPin5 <= slv_reg0(12);
	                   end if;
	               when "PWM"          => 
	                   slv_reg3(17 downto 16) <= "10";
	                   if slv_reg_rden = '1' then
                           if count >= pwmCount then
                                pwmPercent := to_integer(unsigned(slv_reg1(19 downto 16)));
                                pwmCount := 100_000_000/(pwmFrequency5*1000);
                                count := 0;
                           elsif (count <= (pwmCount*pwmPercent/16)) then
                               JAoutputPin5 <= '1';
                           elsif (count > (pwmCount*pwmPercent/16) and (count < (pwmCount))) then
                               JAoutputPin5 <= '0';
                           end if;
	                   end if;
	                   count := count + 1;
	               when "PULSE"        =>
	                   slv_reg3(17 downto 16) <= "01";
	                   if slv_reg_rden = '1' then
	                       if count = 0 then
	                           count := to_integer(unsigned(slv_reg2(19 downto 16)));
	                       end if;
	                       if count > 2 then
	                           JAoutputPin5 <= not JAoutputPin5;
	                       end if;
	                   end if;
	                   if count > 1 then
	                      count := count -1;
	                   end if;
	               when others         =>
	                   slv_reg3(17 downto 16) <= "00";    
	           end case;
	       else 
	           slv_reg3(4) <= '0'; -- busy for JA5
	           count := 0;
	       end if;
	    end if;
	  end if;
	end process;   


	-- JA 6 
	process( S_AXI_ACLK ) is
	variable pwmPercent    : integer := 0;
	variable pwmCount      : integer := 100_000_000/(pwmFrequency6*1000);
	variable count         : integer := 0;
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	       axi_rdata  <= (others => '0');
	    else
	       if slv_reg0(5) = '1' then   -- enable for JA6
	           slv_reg3(5) <= '1';     -- busy for JA6
	           case outType6 is 
	               when "StandardIO"   => 
	                   slv_reg3(19 downto 18) <= "11";
	                   if slv_reg_rden = '1' then
	                       JAoutputPin6 <= slv_reg0(13);
	                   end if;
	               when "PWM"          => 
	                   slv_reg3(19 downto 18) <= "10";
	                   if slv_reg_rden = '1' then
                           if count >= pwmCount then
                                pwmPercent := to_integer(unsigned(slv_reg1(23 downto 20)));
                                pwmCount := 100_000_000/(pwmFrequency6*1000);
                                count := 0;
                           elsif (count <= (pwmCount*pwmPercent/16)) then
                               JAoutputPin6 <= '1';
                           elsif (count > (pwmCount*pwmPercent/16) and (count < (pwmCount))) then
                               JAoutputPin6 <= '0';
                           end if;
	                   end if;
	                   count := count + 1;
	               when "PULSE"        =>
	                   slv_reg3(19 downto 18) <= "01";
	                   if slv_reg_rden = '1' then
	                       if count = 0 then
	                           count := to_integer(unsigned(slv_reg2(23 downto 20)));
	                       end if;
	                       if count > 2 then
	                           JAoutputPin6 <= not JAoutputPin6;
	                       end if;
	                   end if;
	                   if count > 1 then
	                      count := count -1;
	                   end if;
	               when others         =>
	                   slv_reg3(19 downto 18) <= "00";    
	           end case;
	       else 
	           slv_reg3(5) <= '0'; -- busy for JA6
	           count := 0;
	       end if;
	    end if;
	  end if;
	end process;   



	-- JA 7
	process( S_AXI_ACLK ) is
	variable pwmPercent    : integer := 0;
	variable pwmCount      : integer := 100_000_000/(pwmFrequency7*1000);
	variable count         : integer := 0;
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	       axi_rdata  <= (others => '0');
	    else
	       if slv_reg0(6) = '1' then   -- enable for JA7
	           slv_reg3(6) <= '1';     -- busy for JA7
	           case outType7 is 
	               when "StandardIO"   => 
	                   slv_reg3(21 downto 20) <= "11";
	                   if slv_reg_rden = '1' then
	                       JAoutputPin7 <= slv_reg0(14);
	                   end if;
	               when "PWM"          => 
	                   slv_reg3(21 downto 20) <= "10";
	                   if slv_reg_rden = '1' then
                           if count >= pwmCount then
                                pwmPercent := to_integer(unsigned(slv_reg1(29 downto 24)));
                                pwmCount := 100_000_000/(pwmFrequency7*1000);
                                count := 0;
                           elsif (count <= (pwmCount*pwmPercent/16)) then
                               JAoutputPin7 <= '1';
                           elsif (count > (pwmCount*pwmPercent/16) and (count < (pwmCount))) then
                               JAoutputPin7 <= '0';
                           end if;
	                   end if;
	                   count := count + 1;
	               when "PULSE"        =>
	                   slv_reg3(21 downto 20) <= "01";
	                   if slv_reg_rden = '1' then
	                       if count = 0 then
	                           count := to_integer(unsigned(slv_reg2(29 downto 24)));
	                       end if;
	                       if count > 2 then
	                           JAoutputPin7 <= not JAoutputPin7;
	                       end if;
	                   end if;
	                   if count > 1 then
	                      count := count -1;
	                   end if;
	               when others         =>
	                   slv_reg3(21 downto 20) <= "00";    
	           end case;
	       else 
	           slv_reg3(6) <= '0'; -- busy for JA1
	           count := 0;
	       end if;
	    end if;
	  end if;
	end process;   


	-- JA 8
	process( S_AXI_ACLK ) is
	variable pwmPercent    : integer := 0;
	variable pwmCount      : integer := 100_000_000/(pwmFrequency8*1000);
	variable count         : integer := 0;
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	       axi_rdata  <= (others => '0');
	    else
	       if slv_reg0(7) = '1' then   -- enable for JA8
	           slv_reg3(7) <= '1';     -- busy for JA8
	           case outType8 is 
	               when "StandardIO"   => 
	                   slv_reg3(23 downto 22) <= "11";
	                   if slv_reg_rden = '1' then
	                       JAoutputPin8 <= slv_reg0(15);
	                   end if;
	               when "PWM"          => 
	                   slv_reg3(23 downto 22) <= "10";
	                   if slv_reg_rden = '1' then
                           if count >= pwmCount then
                                pwmPercent := to_integer(unsigned(slv_reg1(31 downto 28)));
                                pwmCount := 100_000_000/(pwmFrequency8*1000);
                                count := 0;
                           elsif (count <= (pwmCount*pwmPercent/16)) then
                               JAoutputPin8 <= '1';
                           elsif (count > (pwmCount*pwmPercent/16) and (count < (pwmCount))) then
                               JAoutputPin8 <= '0';
                           end if;
	                   end if;
	                   count := count + 1;
	               when "PULSE"        =>
	                   slv_reg3(23 downto 22) <= "01";
	                   if slv_reg_rden = '1' then
	                       if count = 0 then
	                           count := to_integer(unsigned(slv_reg2(31 downto 28)));
	                       end if;
	                       if count > 2 then
	                           JAoutputPin8 <= not JAoutputPin8;
	                       end if;
	                   end if;
	                   if count > 1 then
	                      count := count -1;
	                   end if;
	               when others         =>
	                   slv_reg3(23 downto 22) <= "00";    
	           end case;
	       else 
	           slv_reg3(7) <= '0'; -- busy for JA1
	           count := 0;
	       end if;
	    end if;
	  end if;
	end process;   



	-- User logic ends

end arch_imp;
